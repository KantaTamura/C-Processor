library IEEE;
use IEEE.std_logic_1164.all;

entity TestALU16 is
end TestALU16;

architecture behavior of TestALU16 is
    constant STEP : Time := 100 ns;

    signal In_A    : std_logic_vector(7 downto 0);
    signal In_B    : std_logic_vector(7 downto 0);
    signal In_C    : std_logic_vector(7 downto 0);
    signal Cin     : std_logic;
    signal modeALU : std_logic_vector(3 downto 0);
    signal Out_F   : std_logic_vector(7 downto 0);
    signal Out_C   : std_logic;
    signal Out_Z   : std_logic;

    component ALU16
        port (
            a    : in  std_logic_vector(7 downto 0);
            b    : in  std_logic_vector(7 downto 0);
            c    : in  std_logic_vector(7 downto 0);
            cin  : in  std_logic;
            mode : in  std_logic_vector(3 downto 0);
            fout : out std_logic_vector(7 downto 0);
            cout : out std_logic;
            zout : out std_logic
        );
    end component;

begin
    ALU : ALU16 port map (In_A, In_B, In_C, Cin, modeALU, Out_F, Out_C, Out_Z);

    process
    begin
        In_A <= "11110000";
        In_B <= "00001111";
        Cin  <= '0';
        modeALU <= "0000";
        wait for STEP;
        modeALU <= "0001";
        wait for STEP;
        modeALU <= "0010";
        wait for STEP;
        modeALU <= "0011";
        wait for STEP;
        modeALU <= "0100";
        wait for STEP;
        modeALU <= "0101";
        wait for STEP;
        modeALU <= "0110";
        wait for STEP;
        modeALU <= "0111";
        wait for STEP;
        modeALU <= "1100";
        wait for STEP;
        modeALU <= "1101";
        wait for STEP;
        modeALU <= "1110";
        wait for STEP;
        modeALU <= "1111";
        wait for STEP;
        modeALU <= "1000";
        wait for STEP;
        modeALU <= "1001";
        wait for STEP;
        modeALU <= "1010";
        wait for STEP;
        modeALU <= "1011";
        wait for STEP;
        In_A    <= "00000010";
        In_B    <= "00000011";
        modeALU <= "0000";
        wait for STEP;
        modeALU <= "0001";
        wait for STEP;
        modeALU <= "0010";
        wait for STEP;
        modeALU <= "0011";
        wait for STEP;
        modeALU <= "0100";
        wait for STEP;
        modeALU <= "0101";
        wait for STEP;
        modeALU <= "0110";
        wait for STEP;
        modeALU <= "0111";
        wait for STEP;
        modeALU <= "1100";
        wait for STEP;
        modeALU <= "1101";
        wait for STEP;
        modeALU <= "1110";
        wait for STEP;
        modeALU <= "1111";
        wait for STEP;
        modeALU <= "1000";
        wait for STEP;
        modeALU <= "1001";
        wait for STEP;
        modeALU <= "1010";
        wait for STEP;
        modeALU <= "1011";
        wait for STEP;
        In_A    <= "00000010";
        In_B    <= "00000011";
        In_C    <= "00000001";
        modeALU <= "1011";
        wait for STEP;
        In_C    <= "00000100";
        modeALU <= "0111";
        wait for STEP;
    wait;
    end process;
end behavior;